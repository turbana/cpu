/* 74283 4-bit adder
 * worse case delay of 80ns
 */
`timescale 1 ns / 100 ps
module \74283 (\1 , \2 , \3 , \4 , \5 , \6 , \7 , \8 , \9 , \10 , \11 , \12 , \13 , \14 , \15 , \16 );
   input \2 , \3  , \5 , \6 , \7 , \8 , \11 , \12 , \14 , \15 , \16 ;
   output \1 , \4 , \9 , \10 , \13 ;

   assign #80 { \9 , \10 , \13 , \1 , \4 } = { 1'b0 , \12 , \14 , \3 , \5 } + { 1'b0 , \11 , \15 , \2 , \6 } + { 1'b0 , 1'b0 , 1'b0 , 1'b0 , \7 };

endmodule
